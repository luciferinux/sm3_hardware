//address decode
module ADDR_DECODER(ENABLE,AHB_HSEL,AHB_HWRITE,REG_ADDR);
output [12:0] ENABLE;
input         AHB_HSEL,AHB_HWRITE;
input  [3:0]  REG_ADDR;
assign ENABLE[0]=AHB_HSEL&AHB_HWRITE&~REG_ADDR[3]&~REG_ADDR[2]&~REG_ADDR[1]&~REG_ADDR[0];
assign ENABLE[1]=AHB_HSEL&AHB_HWRITE&~REG_ADDR[3]&~REG_ADDR[2]&~REG_ADDR[1]&REG_ADDR[0];
assign ENABLE[2]=AHB_HSEL&AHB_HWRITE&~REG_ADDR[3]&~REG_ADDR[2]&REG_ADDR[1]&~REG_ADDR[0];
assign ENABLE[3]=AHB_HSEL&AHB_HWRITE&~REG_ADDR[3]&~REG_ADDR[2]&REG_ADDR[1]&REG_ADDR[0];
assign ENABLE[4]=AHB_HSEL&AHB_HWRITE&~REG_ADDR[3]&REG_ADDR[2]&~REG_ADDR[1]&~REG_ADDR[0];
assign ENABLE[5]=AHB_HSEL&AHB_HWRITE&~REG_ADDR[3]&REG_ADDR[2]&~REG_ADDR[1]&REG_ADDR[0];
assign ENABLE[6]=AHB_HSEL&AHB_HWRITE&~REG_ADDR[3]&REG_ADDR[2]&REG_ADDR[1]&~REG_ADDR[0];
assign ENABLE[7]=AHB_HSEL&AHB_HWRITE&~REG_ADDR[3]&REG_ADDR[2]&REG_ADDR[1]&REG_ADDR[0];
assign ENABLE[8]=AHB_HSEL&AHB_HWRITE&REG_ADDR[3]&~REG_ADDR[2]&~REG_ADDR[1]&~REG_ADDR[0];
assign ENABLE[9]=AHB_HSEL&AHB_HWRITE&REG_ADDR[3]&~REG_ADDR[2]&~REG_ADDR[1]&REG_ADDR[0];
assign ENABLE[10]=AHB_HSEL&AHB_HWRITE&REG_ADDR[3]&~REG_ADDR[2]&REG_ADDR[1]&~REG_ADDR[0];
assign ENABLE[11]=AHB_HSEL&AHB_HWRITE&REG_ADDR[3]&~REG_ADDR[2]&REG_ADDR[1]&REG_ADDR[0];
assign ENABLE[12]=AHB_HSEL&AHB_HWRITE&REG_ADDR[3]&REG_ADDR[2]&~REG_ADDR[1]&~REG_ADDR[0];
endmodule

//REG
module REG(ENABLE,KEY,DAR_ADDR,SAR_ADDR,BSR,CMDR,CRYPT_INTR,AHB_HRDATA,AHB_HRESETN,AHB_HCLK,AHB_HADDR,AHB_HSEL,AHB_HWRITE,SET_STR,AHB_HWDATA);
output          ENABLE,CRYPT_INTR;
output [1:0]    CMDR;
output [12:0]   SAR_ADDR,DAR_ADDR,BSR;
output [31:0]   AHB_HRDATA;
output [191:0]  KEY;
input           AHB_HRESETN,AHB_HCLK,AHB_HSEL,AHB_HWRITE;
input           SET_STR;
input  [5:2]    AHB_HADDR;
input  [31:0]   AHB_HWDATA;
wire            ENR0,STR0,IMR0;
wire   [12:0]   ENABLE_D;
assign CRYPT_INTR=~IMR0&STR0;
assign ENABLE=ENR0;
ADDR_DECODER    addr_decoder(ENABLE_D,AHB_HSEL,AHB_HWRITE,AHB_HADDR);
SDFFldR_1       enr(ENR0,AHB_HWDATA[0],AHB_HCLK,ENABLE_D[0],AHB_HRESETN);
SDFFldR_2       cmdr(CMDR,AHB_HWDATA[1:0],AHB_HCLK,ENABLE_D[1],AHB_HRESETN);
SDFFldR_32      key0(KEY[31:0],AHB_HWDATA,AHB_HCLK,ENABLE_D[2],AHB_HRESETN);
SDFFldR_32      key1(KEY[63:32],AHB_HWDATA,AHB_HCLK,ENABLE_D[3],AHB_HRESETN);
SDFFldR_32      key2(KEY[95:64],AHB_HWDATA,AHB_HCLK,ENABLE_D[4],AHB_HRESETN);
SDFFldR_32      key3(KEY[127:96],AHB_HWDATA,AHB_HCLK,ENABLE_D[5],AHB_HRESETN);
SDFFldR_32      key4(KEY[159:128],AHB_HWDATA,AHB_HCLK,ENABLE_D[6],AHB_HRESETN);
SDFFldR_32      key5(KEY[191:160],AHB_HWDATA,AHB_HCLK,ENABLE_D[7],AHB_HRESETN);
SDFFldR_13      sar(SAR_ADDR,AHB_HWDATA[12:0],AHB_HCLK,ENABLE_D[8],AHB_HRESETN);
SDFFldR_13      dar(DAR_ADDR,AHB_HWDATA[12:0],AHB_HCLK,ENABLE_D[9],AHB_HRESETN);
SDFFldR_13      bsr(BSR,AHB_HWDATA[12:0],AHB_HCLK,ENABLE_D[10],AHB_HRESETN);
SDFFldR_1       str(STR0,SET_STR,AHB_HCLK,ENABLE_D[11],AHB_HRESETN);
SDFFldR_1       imr(IMR0,STR0,AHB_HCLK,ENABLE_D[12],AHB_HRESETN);
MUX1313_32      mux1313_32(AHB_HRDATA,ENR0,CMDR,KEY[31:0],KEY[63:32],KEY[95:64],KEY[127:96],KEY[159:128],KEY[191:160],SAR_ADDR,DAR_ADDR,BSR,IMR0,STR0,ENABLE_D);
endmodule


  


